`timescale 1ns / 1ps 
`include "Procesador_RISC_V.sv"
module test_RISC_V #(Bits = 64, MemSize = 16, N = 32, NumInst = 6); 
  // Inputs
  reg clk, rst; 
  // Creación de una instancia de la unidad bajo prueba (UUT)
  Procesador_RISC_V #(.Bits(Bits), .N(N), .MemSize(MemSize), .NumInst(NumInst)) uut
  (.clk(clk), .rst(rst)); 
  initial 
    begin
      clk = 0;
      $dumpfile("RISCV.vcd");
      $dumpvars(5,uut);
      rst = 0;
      #10
      rst = 1'b1;
      #10
      rst = 1'b0;
      #200
      $finish; 
    end
  always 
    begin
     #5 clk = ~clk; 
    end
    always @(posedge clk) begin 
      prueba(); 
    end 
    task prueba();
	 $monitor("El valor en el registro:")
endmodule

